module register(
	input [15:0] data_in,
	output [15:0] data_out);
