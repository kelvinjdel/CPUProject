module ALU(
	input [15:0] 
